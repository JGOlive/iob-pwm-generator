   // PWM
