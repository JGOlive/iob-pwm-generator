// PWM
output pwm_output
