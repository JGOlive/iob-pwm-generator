   // GPIO
   input [4:0] pwm_input,
   output [4:0] pwm_output,
