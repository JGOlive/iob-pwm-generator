   // PWM

